///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing all MUXs, same 32 inputs
reg[31:0] I[31:0];
wire[31:0] Y2;
wire[31:0] Y3;
wire[31:0] Y4;
wire[31:0] Y8;
wire[31:0] Y32;
reg S2;
reg[1:0] S3;
reg[1:0] S4;
reg[2:0] S8;
reg[4:0] S32;

MUX2_32 myMUX2(.A(I[0]), .B(I[1]), .Y(Y2), .S(S2));
MUX3_32 myMUX3(.A(I[0]), .B(I[1]), .C(I[2]), .Y(Y3), .S(S3));
MUX4_32 myMUX4(.A(I[0]), .B(I[1]), .C(I[2]), .D(I[3]), .Y(Y4), .S(S4));
MUX8_32 myMUX8(.A(I[0]), .B(I[1]), .C(I[2]), .D(I[3]), .E(I[4]), .F(I[5]), .G(I[6]), .H(I[7]), .Y(Y8), .S(S8));
MUX32_32 myMUX32(.I0(I[0]),.I1(I[1]),.I2(I[2]),.I3(I[3]),.I4(I[4]),.I5(I[5]),.I6(I[6]),.I7(I[7]),
.I8(I[8]),.I9(I[9]),.I_10(I[10]),.I_11(I[11]),.I_12(I[12]),.I_13(I[13]),.I_14(I[14]),.I_15(I[15]),
.I_16(I[16]),.I_17(I[17]),.I_18(I[18]),.I_19(I[19]),.I_20(I[20]),.I_21(I[21]),.I_22(I[22]),.I_23(I[23]),
.I_24(I[24]),.I_25(I[25]),.I_26(I[26]),.I_27(I[27]),.I_28(I[28]),.I_29(I[29]),.I_30(I[30]),.I_31(I[31]),.S(S32),.Y(Y32));
//////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// 
integer j;

initial begin

//////////////////////////////////////////////////////////////////////////////
// Initialize 32 input values
for (j = 0; j <= 31; j = j + 1) begin
  I[j] = (2**j)-1;
end
//////////////////////////////////////////////////////////////////////////////

S2 = 1'b1;
S3 = 2'b01;
S4 = 2'b01;
S8 = 3'b001;
S32 = 5'b00001;

#10;
   $display("Testing MUX2");
verifyEqual32(Y2, I[1]);
   $display("Testing MUX3");
verifyEqual32(Y3, I[1]);
   $display("Testing MUX4");
verifyEqual32(Y4, I[1]);
   $display("Testing MUX8");
verifyEqual32(Y8, I[1]);
   $display("Testing MUX32");
verifyEqual32(Y32, I[1]);

 
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule